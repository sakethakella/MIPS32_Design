module execution ();
    
endmodule