module instruction_decode ();
    
endmodule