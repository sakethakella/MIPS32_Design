module memory_access ();
    
endmodule